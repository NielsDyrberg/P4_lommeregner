library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.all;

entity top is
	port(

		clk											: in std_logic
	);

end top;

architecture rtl of top is
	


begin


	
end rtl;




